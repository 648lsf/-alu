module no(out,x);
output [31:0] out;
input [31:0] x;
not not1[31:0](out,x);
// not (out[0],x[0]);
// not (out[1],x[1]);
// not (out[2],x[2]);
// not (out[3],x[3]);
// not (out[4],x[4]);
// not (out[5],x[5]);
// not (out[6],x[6]);
// not (out[7],x[7]);
// not (out[8],x[8]);
// not (out[9],x[9]);
// not (out[10],x[10]);
// not (out[11],x[11]);
// not (out[12],x[12]);
// not (out[13],x[13]);
// not (out[14],x[14]);
// not (out[15],x[15]);
// not (out[16],x[16]);
// not (out[17],x[17]);
// not (out[18],x[18]);
// not (out[19],x[19]);
// not (out[20],x[20]);
// not (out[21],x[21]);
// not (out[22],x[22]);
// not (out[23],x[23]);
// not (out[24],x[24]);
// not (out[25],x[25]);
// not (out[26],x[26]);
// not (out[27],x[27]);
// not (out[28],x[28]);
// not (out[29],x[29]);
// not (out[30],x[30]);
// not (out[31],x[31]);





endmodule